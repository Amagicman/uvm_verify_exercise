`ifndef GPIO_INT_CASE__SV
`define GPIO_INT_CASE__SV

`include "test_gpio_int_int_code.sv"
`include "test_gpio_int_reg_rw.sv"
`include "test_gpio_int_priority.sv"
`include "test_gpio_int_oriented.sv"

`endif

`ifndef GPIO_INT_CASE__SV
`define GPIO_INT_CASE__SV

`include "test_reg_rw.sv"
`include "test_intr_code.sv"
`include "test_int_same_domain_multi.sv"
`include "test_int_same_cont.sv"
`include "test_gpio_int_cov.sv"
`include "test_int_priority.sv"

`endif
